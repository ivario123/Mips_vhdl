library IEEE;
use IEEE.std_logic_1164.all;

entity programmemory is
  port( address:in std_logic_vector(31 downto 0);
        instruction: out std_logic_vector(31 downto 0)
        );
end programmemory;

architecture behav of programmemory is
begin

with address select
-- Base test
      instruction <=    "00100000001000001111111111111000" when X"00000000", --addi r0,r1,-8
                        "00100000010000010000000000000011" when X"00000004", --addi r1,r2,3
                        "00000000000000010001000000100000" when X"00000008", --add r2,r0,r1
                        "00000000001000000001100000100010" when X"0000000c", --sub r3,r1,r0
                        "00000000010000110010000000101010" when X"00000010", --slt r4,r2,r3
                        "00101000010001001111111111110111" when X"00000014", --slti r4,r2,-9
                        "00000000010000110010000000101010" when X"00000018", --slt r4,r2,r3
                        "00000000100001100010100000100101" when X"0000001c", --or  r5,r4,r6
                        "00000000101000010011000000100100" when X"00000020", --and r6,r5,r1
                        "10101100111000100000000000000000" when X"00000024", -- sw r2, 0(r7) 
                        "10001100111010000000000000000000" when X"00000028", -- lw r8, 0(r7)  
                        "10101101001000110000000000000100" when X"0000002c", -- sw r3, 4(r9)
                        "10001101010010010000000000000100" when X"00000030", -- lw r9, 4(r10)
                        "11111100001000000000000000000001" when others;
    
--    instruction <=  -- N =  12 and D =  5  to change what 2 numbers are devided change the X"00000000" and X"00000004" instructions
--                    "00100000000001000000000000001100" when X"00000000", -- addi $a0, $0, N; addi $t, $s, imm   
--                    "00100000000001010000000000000101" when X"00000004", -- addi $a1, $0, D; addi $t, $s, imm     
--                    -- N = 12 D = 12
--                    --"00100000000001000000000000001100" when X"00000000", -- addi $a0, $0, N; addi $t, $s, imm   
--                    --"00100000000001010000000000001100" when X"00000004", -- addi $a1, $0, D; addi $t, $s, imm   
--                    -- N = 5 and D = 12
--                    --"00100000000001000000000000000101" when X"00000000", -- addi $a0, $0, N; addi $t, $s, imm   
--                    --"00100000000001010000000000001100" when X"00000004", -- addi $a1, $0, D; addi $t, $s, imm   
--                    -- Do not comment out
--                    "00100000000001100000000000000001" when X"00000008", -- addi $a2, $0, 0x0001; addi $t, $s, imm     
--                    "00000000000000000001000000100000" when X"0000000c",  -- add $v0, $0, $0; add $d, $s, $t   
--                    "00000000000001000001100000100000" when X"00000010", -- add $v1, $0, $a0; add $d, $s, $t   
--                    "00000000011001010100000000101010" when X"00000014", -- slt $t0, $v1, $a0;slt $d, $s, $t
--                    "00010001000001100000000000000100" when X"00000018", -- beq $t0, $a2, 0x0005;beq $s, $t, offset  
--                    "00100000010000100000000000000001" when X"0000001c", -- addi $v0, $v0, 0x0001; addi $t, $s, imm       
--                    "00000000011001010001100000100010" when X"00000020", -- sub $v1, $v1, $a1; sub $d, $s, $t  
--                    "00001000000000000000000000000101" when X"00000024", -- J 6
--                    "00000000000000000000000000000000" when others; -- Noop
    
   
                            
end behav;